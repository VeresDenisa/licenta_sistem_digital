package CS_environment_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import item_pack::*;
    import CS_sequence_pack::*;

    import CS_agent_pack::*;
    import CS_coverage_pack::*;
    
    `include "testbench/CS/test/environment/CS_environment.svh"

  endpackage : CS_environment_pack
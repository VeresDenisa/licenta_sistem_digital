package LM_environment_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import item_pack::*;
    import LM_sequence_pack::*;
  
    import LM_agent_pack::*;
    import LM_coverage_pack::*;
   
    `include "testbench/environment_config.svh"

    `include "testbench/LM/test/environment/LM_environment.svh"
  endpackage : LM_environment_pack
package UART_coverage_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import item_pack::*;
  
    `include "testbench/UART/test/environment/coverage/UART_covergroup.sv"
    
    `include "testbench/UART/test/environment/coverage/UART_coverage.svh"
  endpackage : UART_coverage_pack
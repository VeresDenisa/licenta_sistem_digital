package DB_agent_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import item_pack::*;
  
    `include "testbench/agent_config.svh"

    `include "testbench/DB/test/environment/agent/DB_driver.svh"
    `include "testbench/DB/test/environment/agent/DB_monitor.svh"
    `include "testbench/DB/test/environment/agent/DB_agent.svh"
  endpackage : DB_agent_pack










package CD_sequence_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import item_pack::*;
  
    `include "testbench/CM/test/sequence/CM_input_sequence.svh"

    `include "testbench/CONF/test/sequence/CONF_input_sequence.svh"
  endpackage : CD_sequence_pack
package DB_coverage_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import item_pack::*;
  
    `include "testbench/DB/test/environment/coverage/DB_covergroup.sv"

    `include "testbench/DB/test/environment/coverage/DB_coverage.svh"
  endpackage : DB_coverage_pack
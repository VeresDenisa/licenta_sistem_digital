package LM_sequence_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import item_pack::*;
  
    `include "testbench/CM/test/sequence/CM_output_sequence.svh"

    `include "testbench/UART/test/sequence/UART_output_sequence.svh"
  endpackage : LM_sequence_pack
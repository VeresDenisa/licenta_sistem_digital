package VGA_coverage_pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    import item_pack::*;
  
    `include "testbench/VGA/test/environment/coverage/VGA_covergroup.sv"

    `include "testbench/VGA/test/environment/coverage/VGA_coverage.svh"
  endpackage : VGA_coverage_pack